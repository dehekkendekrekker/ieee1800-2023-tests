module miter (
  input  [  0:0] \__pi_dummy ,
`ifdef DIRECT_CROSS_POINTS
`else
`endif
  output [  0:0] \__mp_a__gold ,
  output [  0:0] \__mp_a__gate
);
  \gold.simple_immediate_assert_statement gold (
    .\__pi_dummy (\__pi_dummy ),
`ifdef DIRECT_CROSS_POINTS
`else
`endif
    .\__mp_a (\__mp_a__gold )
  );
  \gate.simple_immediate_assert_statement gate (
    .\__pi_dummy (\__pi_dummy ),
`ifdef DIRECT_CROSS_POINTS
`else
`endif
    .\__mp_a (\__mp_a__gate )
  );
`ifdef ASSUME_DEFINED_INPUTS
  miter_def_prop #(1, "assume") \__pi_dummy__assume (\__pi_dummy );
`endif
`ifndef DIRECT_CROSS_POINTS
`endif
`ifdef CHECK_MATCH_POINTS
  miter_cmp_prop #(1, "assert") \__mp_a__assert (\__mp_a__gold , \__mp_a__gate );
`endif
`ifdef CHECK_OUTPUTS
`endif
`ifdef COVER_DEF_CROSS_POINTS
  `ifdef DIRECT_CROSS_POINTS
  `else
  `endif
`endif
`ifdef COVER_DEF_GOLD_MATCH_POINTS
  miter_def_prop #(1, "cover") \__mp_a__gold_cover (\__mp_a__gold );
`endif
`ifdef COVER_DEF_GATE_MATCH_POINTS
  miter_def_prop #(1, "cover") \__mp_a__gate_cover (\__mp_a__gate );
`endif
`ifdef COVER_DEF_GOLD_OUTPUTS
`endif
`ifdef COVER_DEF_GATE_OUTPUTS
`endif
endmodule
module miter_cmp_prop #(parameter WIDTH=1, parameter TYPE="assert") (input [WIDTH-1:0] in_gold, in_gate);
  reg okay;
  integer i;
  always @* begin
    okay = 1;
    for (i = 0; i < WIDTH; i = i+1)
      okay = okay && (in_gold[i] === 1'bx || in_gold[i] === in_gate[i]);
  end
  generate
    if (TYPE == "assert") always @* assert(okay);
    if (TYPE == "assume") always @* assume(okay);
    if (TYPE == "cover")  always @* cover(okay);
  endgenerate
endmodule
module miter_def_prop #(parameter WIDTH=1, parameter TYPE="assert") (input [WIDTH-1:0] in);
  wire okay = ^in !== 1'bx;
  generate
    if (TYPE == "assert") always @* assert(okay);
    if (TYPE == "assume") always @* assume(okay);
    if (TYPE == "cover")  always @* cover(okay);
  endgenerate
endmodule
module \gold.simple_immediate_assert_statement (
  input  [  0:0] \__pi_dummy ,
  output [  0:0] \__mp_a
);
endmodule
module \gate.simple_immediate_assert_statement (
  input  [  0:0] \__pi_dummy ,
  output [  0:0] \__mp_a
);
endmodule
